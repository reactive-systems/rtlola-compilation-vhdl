library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.fixed_pkg.all;
use work.array_type_pkg.all;

entity queue is
    port (
        clk, rst : in std_logic;
        push : in std_logic;
        time_data_in : in unsigned(63 downto 0);
		a_data_in : in std_logic;
		a_en_in : in std_logic;
		b_data_in : in std_logic;
		b_en_in : in std_logic;
		ID_data_in : in signed(7 downto 0);
		ID_en_in : in std_logic;
		eq_en_in : in std_logic;
		lt_en_in : in std_logic;
		le_en_in : in std_logic;
		gt_en_in : in std_logic;
		ge_en_in : in std_logic;
		neq_en_in : in std_logic;
		not_a_en_in : in std_logic;
		a_and_b_en_in : in std_logic;
		a_or_b_en_in : in std_logic;
		a_impl_b_en_in : in std_logic;
		a_equiv_b_en_in : in std_logic;
		a_xor_b_en_in : in std_logic;
		true_const_en_in : in std_logic;
		time_stream_en_in : in std_logic;
        full : out std_logic;
        pop : in std_logic;
        time_data_out : out unsigned(63 downto 0);
		a_data_out : out std_logic;
		a_en_out : out std_logic;
		b_data_out : out std_logic;
		b_en_out : out std_logic;
		ID_data_out : out signed(7 downto 0);
		ID_en_out : out std_logic;
		eq_en_out : out std_logic;
		lt_en_out : out std_logic;
		le_en_out : out std_logic;
		gt_en_out : out std_logic;
		ge_en_out : out std_logic;
		neq_en_out : out std_logic;
		not_a_en_out : out std_logic;
		a_and_b_en_out : out std_logic;
		a_or_b_en_out : out std_logic;
		a_impl_b_en_out : out std_logic;
		a_equiv_b_en_out : out std_logic;
		a_xor_b_en_out : out std_logic;
		true_const_en_out : out std_logic;
		time_stream_en_out : out std_logic;
        available : out std_logic
    );
end queue;

architecture behavioral of queue is

    signal is_full : std_logic;
    signal time_data_reg : unsigned64_array(1 downto 0);
    signal time_data : unsigned(63 downto 0);
	signal a_data_reg : bit_array(1 downto 0);
	signal a_en_reg : bit_array(1 downto 0);
	signal a_data : std_logic;
	signal a_en: std_logic;
	signal b_data_reg : bit_array(1 downto 0);
	signal b_en_reg : bit_array(1 downto 0);
	signal b_data : std_logic;
	signal b_en: std_logic;
	signal ID_data_reg : signed8_array(1 downto 0);
	signal ID_en_reg : bit_array(1 downto 0);
	signal ID_data : signed(7 downto 0);
	signal ID_en: std_logic;
	signal eq_en_reg : bit_array(1 downto 0);
	signal eq_en : std_logic;
	signal lt_en_reg : bit_array(1 downto 0);
	signal lt_en : std_logic;
	signal le_en_reg : bit_array(1 downto 0);
	signal le_en : std_logic;
	signal gt_en_reg : bit_array(1 downto 0);
	signal gt_en : std_logic;
	signal ge_en_reg : bit_array(1 downto 0);
	signal ge_en : std_logic;
	signal neq_en_reg : bit_array(1 downto 0);
	signal neq_en : std_logic;
	signal not_a_en_reg : bit_array(1 downto 0);
	signal not_a_en : std_logic;
	signal a_and_b_en_reg : bit_array(1 downto 0);
	signal a_and_b_en : std_logic;
	signal a_or_b_en_reg : bit_array(1 downto 0);
	signal a_or_b_en : std_logic;
	signal a_impl_b_en_reg : bit_array(1 downto 0);
	signal a_impl_b_en : std_logic;
	signal a_equiv_b_en_reg : bit_array(1 downto 0);
	signal a_equiv_b_en : std_logic;
	signal a_xor_b_en_reg : bit_array(1 downto 0);
	signal a_xor_b_en : std_logic;
	signal true_const_en_reg : bit_array(1 downto 0);
	signal true_const_en : std_logic;
	signal time_stream_en_reg : bit_array(1 downto 0);
	signal time_stream_en : std_logic;
    signal av : std_logic;
    signal size : integer;
    signal clk_reg : std_logic;
    signal push_done : std_logic;
    signal pop_done : std_logic;

begin

    process(rst, clk) begin
        if (rst = '1') then
            is_full <= '0';
            time_data_reg(time_data_reg'high downto 0) <= (others => (others => '0'));
            time_data <= (others => '0');
			a_data_reg(a_data_reg'high downto 0) <= (others => '0');
			a_en_reg(a_en_reg'high downto 0) <= (others => '0');
			a_data <= '0';
			a_en <= '0';
			b_data_reg(b_data_reg'high downto 0) <= (others => '0');
			b_en_reg(b_en_reg'high downto 0) <= (others => '0');
			b_data <= '0';
			b_en <= '0';
			ID_data_reg(ID_data_reg'high downto 0) <= (others => (others => '0'));
			ID_en_reg(ID_en_reg'high downto 0) <= (others => '0');
			ID_data <= (others => '0');
			ID_en <= '0';
			eq_en_reg <= (others => '0');
			eq_en <= '0';
			lt_en_reg <= (others => '0');
			lt_en <= '0';
			le_en_reg <= (others => '0');
			le_en <= '0';
			gt_en_reg <= (others => '0');
			gt_en <= '0';
			ge_en_reg <= (others => '0');
			ge_en <= '0';
			neq_en_reg <= (others => '0');
			neq_en <= '0';
			not_a_en_reg <= (others => '0');
			not_a_en <= '0';
			a_and_b_en_reg <= (others => '0');
			a_and_b_en <= '0';
			a_or_b_en_reg <= (others => '0');
			a_or_b_en <= '0';
			a_impl_b_en_reg <= (others => '0');
			a_impl_b_en <= '0';
			a_equiv_b_en_reg <= (others => '0');
			a_equiv_b_en <= '0';
			a_xor_b_en_reg <= (others => '0');
			a_xor_b_en <= '0';
			true_const_en_reg <= (others => '0');
			true_const_en <= '0';
			time_stream_en_reg <= (others => '0');
			time_stream_en <= '0';
            size <= 0;
            av <= '0';
            clk_reg <= '0';
            push_done <= '0';
            pop_done <= '0';
        elsif rising_edge(clk) then
            clk_reg <= not clk_reg;
            if clk_reg = '0' then
                if push = '1' and push_done = '0' and pop = '1' and pop_done = '0' and size > 0 and size < 2 then
                    -- perform push and pop
                    time_data_reg <= time_data_reg(time_data_reg'high - 1 downto 0) & time_data_in;
					a_data_reg <= a_data_reg(a_data_reg'high - 1 downto 0) & a_data_in;
					a_en_reg <= a_en_reg(a_en_reg'high - 1 downto 0) & a_en_in;
					b_data_reg <= b_data_reg(b_data_reg'high - 1 downto 0) & b_data_in;
					b_en_reg <= b_en_reg(b_en_reg'high - 1 downto 0) & b_en_in;
					ID_data_reg <= ID_data_reg(ID_data_reg'high - 1 downto 0) & ID_data_in;
					ID_en_reg <= ID_en_reg(ID_en_reg'high - 1 downto 0) & ID_en_in;
					eq_en_reg <= eq_en_reg(eq_en_reg'high - 1 downto 0) & eq_en_in;
					lt_en_reg <= lt_en_reg(lt_en_reg'high - 1 downto 0) & lt_en_in;
					le_en_reg <= le_en_reg(le_en_reg'high - 1 downto 0) & le_en_in;
					gt_en_reg <= gt_en_reg(gt_en_reg'high - 1 downto 0) & gt_en_in;
					ge_en_reg <= ge_en_reg(ge_en_reg'high - 1 downto 0) & ge_en_in;
					neq_en_reg <= neq_en_reg(neq_en_reg'high - 1 downto 0) & neq_en_in;
					not_a_en_reg <= not_a_en_reg(not_a_en_reg'high - 1 downto 0) & not_a_en_in;
					a_and_b_en_reg <= a_and_b_en_reg(a_and_b_en_reg'high - 1 downto 0) & a_and_b_en_in;
					a_or_b_en_reg <= a_or_b_en_reg(a_or_b_en_reg'high - 1 downto 0) & a_or_b_en_in;
					a_impl_b_en_reg <= a_impl_b_en_reg(a_impl_b_en_reg'high - 1 downto 0) & a_impl_b_en_in;
					a_equiv_b_en_reg <= a_equiv_b_en_reg(a_equiv_b_en_reg'high - 1 downto 0) & a_equiv_b_en_in;
					a_xor_b_en_reg <= a_xor_b_en_reg(a_xor_b_en_reg'high - 1 downto 0) & a_xor_b_en_in;
					true_const_en_reg <= true_const_en_reg(true_const_en_reg'high - 1 downto 0) & true_const_en_in;
					time_stream_en_reg <= time_stream_en_reg(time_stream_en_reg'high - 1 downto 0) & time_stream_en_in;

                    time_data <= time_data_reg(size-1);
					a_data <= a_data_reg(size-1);
					a_en <= a_en_reg(size-1);
					b_data <= b_data_reg(size-1);
					b_en <= b_en_reg(size-1);
					ID_data <= ID_data_reg(size-1);
					ID_en <= ID_en_reg(size-1);
					eq_en <= eq_en_reg(size-1);
					lt_en <= lt_en_reg(size-1);
					le_en <= le_en_reg(size-1);
					gt_en <= gt_en_reg(size-1);
					ge_en <= ge_en_reg(size-1);
					neq_en <= neq_en_reg(size-1);
					not_a_en <= not_a_en_reg(size-1);
					a_and_b_en <= a_and_b_en_reg(size-1);
					a_or_b_en <= a_or_b_en_reg(size-1);
					a_impl_b_en <= a_impl_b_en_reg(size-1);
					a_equiv_b_en <= a_equiv_b_en_reg(size-1);
					a_xor_b_en <= a_xor_b_en_reg(size-1);
					true_const_en <= true_const_en_reg(size-1);
					time_stream_en <= time_stream_en_reg(size-1);
                    push_done <= '1';
                    pop_done <= '1';
                elsif push = '1' and push_done = '0' and size < 2 then
                    -- perform push
                    time_data_reg <= time_data_reg(time_data_reg'high - 1 downto 0) & time_data_in;
					a_data_reg <= a_data_reg(a_data_reg'high - 1 downto 0) & a_data_in;
					a_en_reg <= a_en_reg(a_en_reg'high - 1 downto 0) & a_en_in;
					b_data_reg <= b_data_reg(b_data_reg'high - 1 downto 0) & b_data_in;
					b_en_reg <= b_en_reg(b_en_reg'high - 1 downto 0) & b_en_in;
					ID_data_reg <= ID_data_reg(ID_data_reg'high - 1 downto 0) & ID_data_in;
					ID_en_reg <= ID_en_reg(ID_en_reg'high - 1 downto 0) & ID_en_in;
					eq_en_reg <= eq_en_reg(eq_en_reg'high - 1 downto 0) & eq_en_in;
					lt_en_reg <= lt_en_reg(lt_en_reg'high - 1 downto 0) & lt_en_in;
					le_en_reg <= le_en_reg(le_en_reg'high - 1 downto 0) & le_en_in;
					gt_en_reg <= gt_en_reg(gt_en_reg'high - 1 downto 0) & gt_en_in;
					ge_en_reg <= ge_en_reg(ge_en_reg'high - 1 downto 0) & ge_en_in;
					neq_en_reg <= neq_en_reg(neq_en_reg'high - 1 downto 0) & neq_en_in;
					not_a_en_reg <= not_a_en_reg(not_a_en_reg'high - 1 downto 0) & not_a_en_in;
					a_and_b_en_reg <= a_and_b_en_reg(a_and_b_en_reg'high - 1 downto 0) & a_and_b_en_in;
					a_or_b_en_reg <= a_or_b_en_reg(a_or_b_en_reg'high - 1 downto 0) & a_or_b_en_in;
					a_impl_b_en_reg <= a_impl_b_en_reg(a_impl_b_en_reg'high - 1 downto 0) & a_impl_b_en_in;
					a_equiv_b_en_reg <= a_equiv_b_en_reg(a_equiv_b_en_reg'high - 1 downto 0) & a_equiv_b_en_in;
					a_xor_b_en_reg <= a_xor_b_en_reg(a_xor_b_en_reg'high - 1 downto 0) & a_xor_b_en_in;
					true_const_en_reg <= true_const_en_reg(true_const_en_reg'high - 1 downto 0) & true_const_en_in;
					time_stream_en_reg <= time_stream_en_reg(time_stream_en_reg'high - 1 downto 0) & time_stream_en_in;

                    size <= size + 1;
                    av <= '1';
                    is_full <= to_std_logic(size = 1);
                    push_done <= '1';
                elsif pop = '1' and pop_done = '0' and size > 0 then
                    --perform pop
                    time_data <= time_data_reg(size-1);
					a_data <= a_data_reg(size-1);
					a_en <= a_en_reg(size-1);
					b_data <= b_data_reg(size-1);
					b_en <= b_en_reg(size-1);
					ID_data <= ID_data_reg(size-1);
					ID_en <= ID_en_reg(size-1);
					eq_en <= eq_en_reg(size-1);
					lt_en <= lt_en_reg(size-1);
					le_en <= le_en_reg(size-1);
					gt_en <= gt_en_reg(size-1);
					ge_en <= ge_en_reg(size-1);
					neq_en <= neq_en_reg(size-1);
					not_a_en <= not_a_en_reg(size-1);
					a_and_b_en <= a_and_b_en_reg(size-1);
					a_or_b_en <= a_or_b_en_reg(size-1);
					a_impl_b_en <= a_impl_b_en_reg(size-1);
					a_equiv_b_en <= a_equiv_b_en_reg(size-1);
					a_xor_b_en <= a_xor_b_en_reg(size-1);
					true_const_en <= true_const_en_reg(size-1);
					time_stream_en <= time_stream_en_reg(size-1);

                    size <= size - 1;
                    is_full <= '0';
                    av <= to_std_logic(size > 1);
                    pop_done <= '1';
                end if;
            else
                if push = '0' then
                    push_done <= '0';
                end if;
                if pop = '0' then 
                    pop_done <= '0';
                end if;
            end if;
        end if;
    end process;

    full <= is_full;
    time_data_out <= time_data;
	a_data_out <= a_data;
	a_en_out <= a_en;
	b_data_out <= b_data;
	b_en_out <= b_en;
	ID_data_out <= ID_data;
	ID_en_out <= ID_en;
	eq_en_out <= eq_en;
	lt_en_out <= lt_en;
	le_en_out <= le_en;
	gt_en_out <= gt_en;
	ge_en_out <= ge_en;
	neq_en_out <= neq_en;
	not_a_en_out <= not_a_en;
	a_and_b_en_out <= a_and_b_en;
	a_or_b_en_out <= a_or_b_en;
	a_impl_b_en_out <= a_impl_b_en;
	a_equiv_b_en_out <= a_equiv_b_en;
	a_xor_b_en_out <= a_xor_b_en;
	true_const_en_out <= true_const_en;
	time_stream_en_out <= time_stream_en;
    available <= av;

end behavioral;
